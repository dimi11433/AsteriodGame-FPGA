library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Types.all;

entity get_character_rom is
    port (
        char_addr : in std_logic_vector(7 downto 0);
        char_data : out char_bitmap
    );
end entity get_character_rom;

architecture rom of get_character_rom is
    -- char_bitmap type is now declared in Font_Types package.
    -- Define a type for the complete font ROM: 26 letters + 10 digits = 36 characters.
    type font_rom_type is array (0 to 64) of char_bitmap;

    -- FONT_ROM: array mapping character indices (0-64) to 8x8 bitmap patterns for '0'-'9', 'a'-'z', and 'A'-'Z'
    constant FONT_ROM : font_rom_type := (
        -- '0'
        0 => (
        "00111000",
        "01000100",
        "01001100",
        "01010100",
        "01100100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '1'
        1 => (
        "00010000",
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- '2'
        2 => (
        "00111000",
        "01000100",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "01111100",
        "00000000"
        ),
        -- '3'
        3 => (
        "00111000",
        "01000100",
        "00000100",
        "00011000",
        "00000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '4'
        4 => (
        "00001000",
        "00011000",
        "00101000",
        "01001000",
        "01111100",
        "00001000",
        "00001000",
        "00000000"
        ),
        -- '5'
        5 => (
        "01111100",
        "01000000",
        "01111000",
        "00000100",
        "00000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '6'
        6 => (
        "00111000",
        "01000000",
        "01000000",
        "01111000",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '7'
        7 => (
        "01111100",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "00100000",
        "00100000",
        "00000000"
        ),
        -- '8'
        8 => (
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '9'
        9 => (
        "00111000",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'a'
        10 => (
        "00000000",
        "00000000",
        "00111000",
        "00000100",
        "00111100",
        "01000100",
        "00111100",
        "00000000"
        ),
        -- 'b'
        11 => (
        "01000000",
        "01000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01110000",
        "00000000"
        ),
        -- 'c'
        12 => (
        "00000000",
        "00000000",
        "00111000",
        "01000000",
        "01000000",
        "01000000",
        "00111000",
        "00000000"
        ),
        -- 'd'
        13 => (
        "00000100",
        "00000100",
        "00110100",
        "01001100",
        "01000100",
        "01000100",
        "00111100",
        "00000000"
        ),
        -- 'e'
        14 => (
        "00000000",
        "00000000",
        "00111000",
        "01000100",
        "01111000",
        "01000000",
        "00111000",
        "00000000"
        ),
        -- 'f'
        15 => (
        "00011000",
        "00100000",
        "01110000",
        "00100000",
        "00100000",
        "00100000",
        "00100000",
        "00000000"
        ),
        -- 'g'
        16 => (
        "00000000",
        "00111100",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'h'
        17 => (
        "01000000",
        "01000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00000000"
        ),
        -- 'i'
        18 => (
        "00010000",
        "00000000",
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- 'j'
        19 => (
        "00001000",
        "00000000",
        "00011000",
        "00001000",
        "00001000",
        "01001000",
        "00110000",
        "00000000"
        ),
        -- 'k'
        20 => (
        "01000000",
        "01010000",
        "01100000",
        "01110000",
        "01011000",
        "01001000",
        "01000100",
        "00000000"
        ),
        -- 'l'
        21 => (
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- 'm'
        22 => (
        "00000000",
        "00000000",
        "01101000",
        "01010100",
        "01010100",
        "01010100",
        "01010100",
        "00000000"
        ),
        -- 'n'
        23 => (
        "00000000",
        "00000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00000000"
        ),
        -- 'o'
        24 => (
        "00000000",
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- 'p'
        25 => (
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "01000000",
        "01000000",
        "00000000"
        ),
        -- 'q'
        26 => (
        "00000000",
        "00111100",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00000000"
        ),
        -- 'r'
        27 => (
        "00000000",
        "00000000",
        "01011000",
        "01100100",
        "01000000",
        "01000000",
        "01000000",
        "00000000"
        ),
        -- 's'
        28 => (
        "00000000",
        "00000000",
        "00111100",
        "01000000",
        "00111000",
        "00000100",
        "01111000",
        "00000000"
        ),
        -- 't'
        29 => (
        "00100000",
        "00100000",
        "01110000",
        "00100000",
        "00100000",
        "00100000",
        "00011000",
        "00000000"
        ),
        -- 'u'
        30 => (
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00111000",
        "00000000"
        ),
        -- 'v'
        31 => (
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "01001000",
        "00110000",
        "00010000",
        "00000000"
        ),
        -- 'w'
        32 => (
        "00000000",
        "00000000",
        "01000100",
        "01010100",
        "01010100",
        "01111100",
        "01000100",
        "00000000"
        ),
        -- 'x'
        33 => (
        "00000000",
        "00000000",
        "01000100",
        "00101000",
        "00010000",
        "00101000",
        "01000100",
        "00000000"
        ),
        -- 'y'
        34 => (
        "00000000",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'z'
        35 => (
        "00000000",
        "00000000",
        "01111100",
        "00001000",
        "00010000",
        "00100000",
        "01111100",
        "00000000"
        ),
        -- 'A'
        36 => (
            "00011000",
            "00100100",
            "01000010",
            "01000010",
            "01111110",
            "01000010",
            "01000010",
            "00000000"
        ),
        -- 'B'
        37 => (
            "01111000",
            "01000100",
            "01000100",
            "01111000",
            "01000100",
            "01000100",
            "01111000",
            "00000000"
        ),
        -- 'C'
        38 => (
            "00111100",
            "01000010",
            "01000000",
            "01000000",
            "01000000",
            "01000010",
            "00111100",
            "00000000"
        ),
        -- 'D'
        39 => (
            "01111000",
            "01000100",
            "01000010",
            "01000010",
            "01000010",
            "01000100",
            "01111000",
            "00000000"
        ),
        -- 'E'
        40 => (
            "01111110",
            "01000000",
            "01000000",
            "01111100",
            "01000000",
            "01000000",
            "01111110",
            "00000000"
        ),
        -- 'F'
        41 => (
            "01111110",
            "01000000",
            "01000000",
            "01111100",
            "01000000",
            "01000000",
            "01000000",
            "00000000"
        ),
        -- 'G'
        42 => (
            "00111100",
            "01000010",
            "01000000",
            "01001110",
            "01000010",
            "01000010",
            "00111100",
            "00000000"
        ),
        -- 'H'
        43 => (
            "01000010",
            "01000010",
            "01000010",
            "01111110",
            "01000010",
            "01000010",
            "01000010",
            "00000000"
        ),
        -- 'I'
        44 => (
            "00111000",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00111000",
            "00000000"
        ),
        -- 'J'
        45 => (
            "00011110",
            "00000100",
            "00000100",
            "00000100",
            "01000100",
            "01000100",
            "00111000",
            "00000000"
        ),
        -- 'K'
        46 => (
            "01000010",
            "01000100",
            "01001000",
            "01110000",
            "01001000",
            "01000100",
            "01000010",
            "00000000"
        ),
        -- 'L'
        47 => (
            "01000000",
            "01000000",
            "01000000",
            "01000000",
            "01000000",
            "01000000",
            "01111110",
            "00000000"
        ),
        -- 'M'
        48 => (
            "01000010",
            "01100110",
            "01011010",
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "00000000"
        ),
        -- 'N'
        49 => (
            "01000010",
            "01100010",
            "01010010",
            "01001010",
            "01000110",
            "01000010",
            "01000010",
            "00000000"
        ),
        -- 'O'
        50 => (
            "00111100",
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "00111100",
            "00000000"
        ),
        -- 'P'
        51 => (
            "01111100",
            "01000010",
            "01000010",
            "01111100",
            "01000000",
            "01000000",
            "01000000",
            "00000000"
        ),
        -- 'Q'
        52 => (
            "00111100",
            "01000010",
            "01000010",
            "01000010",
            "01001010",
            "00111100",
            "00000010",
            "00000000"
        ),
        -- 'R'
        53 => (
            "01111100",
            "01000010",
            "01000010",
            "01111100",
            "01001000",
            "01000100",
            "01000010",
            "00000000"
        ),
        -- 'S'
        54 => (
            "00111100",
            "01000010",
            "01000000",
            "00111100",
            "00000010",
            "01000010",
            "00111100",
            "00000000"
        ),
        -- 'T'
        55 => (
            "01111110",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00000000"
        ),
        -- 'U'
        56 => (
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "00111100",
            "00000000"
        ),
        -- 'V'
        57 => (
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "01000010",
            "00100100",
            "00011000",
            "00000000"
        ),
        -- 'W'
        58 => (
            "01000010",
            "01000010",
            "01000010",
            "01011010",
            "01011010",
            "01100110",
            "01000010",
            "00000000"
        ),
        -- 'X'
        59 => (
            "01000010",
            "00100100",
            "00011000",
            "00011000",
            "00011000",
            "00100100",
            "01000010",
            "00000000"
        ),
        -- 'Y'
        60 => (
            "01000010",
            "00100100",
            "00011000",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00000000"
        ),
        -- 'Z'
        61 => (
            "01111110",
            "00000100",
            "00001000",
            "00010000",
            "00100000",
            "01000000",
            "01111110",
            "00000000"
        ),
        -- ',' (comma)
        62 => (
            "00000000",
            "00000000",
            "00000000",
            "00000000",
            "00000000",
            "00010000",
            "00010000",
            "00100000"
        ),
        -- '.' (period)
        63 => (
            "00000000",
            "00000000",
            "00000000",
            "00000000",
            "00000000",
            "00000000",
            "00110000",
            "00110000"
        ),
        -- '!' (exclamation)
        64 => (
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00010000",
            "00000000",
            "00010000",
            "00000000"
        )
    );
    -- Convert 8-bit char_addr to integer index for ROM lookup
    signal index : integer;
begin
    -- Compute ROM index from input address vector
    index <= to_integer(unsigned(char_addr));

    -- Process to index into FONT_ROM using char_addr
    -- ROM access process: select bitmap based on computed index
    process (index)
    begin
        -- Range check: if index is within valid ROM entries
        if index < 65 and index >= 0 then
            -- Assign corresponding character bitmap from ROM
            char_data <= FONT_ROM(index);
        -- If index is out of range, output blank bitmap (all zeros)
        else
            char_data <= (others => (others => '0'));
        end if;
    end process;

end rom;