-- Package Declaration
package Font_Types is
    type char_bitmap is array (0 to 7) of std_logic_vector(7 downto 0);
end package Font_Types;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity get_character_rom is
    port (
        char_addr : in std_logic_vector(7 downto 0);
        char_data : out char_bitmap
    );
end entity get_character_rom;

architecture rom of get_character_rom is
    -- char_bitmap type is now declared in Font_Types package.
    -- Define a type for the complete font ROM: 26 letters + 10 digits = 36 characters.
    type font_rom_type is array (0 to 35) of char_bitmap;

    constant FONT_ROM : font_rom_type := (
        -- 'a'
        0 => (
        "00000000",
        "00000000",
        "00111000",
        "00000100",
        "00111100",
        "01000100",
        "00111100",
        "00000000"
        ),
        -- 'b'
        1 => (
        "01000000",
        "01000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01110000",
        "00000000"
        ),
        -- 'c'
        2 => (
        "00000000",
        "00000000",
        "00111000",
        "01000000",
        "01000000",
        "01000000",
        "00111000",
        "00000000"
        ),
        -- 'd'
        3 => (
        "00000100",
        "00000100",
        "00110100",
        "01001100",
        "01000100",
        "01000100",
        "00111100",
        "00000000"
        ),
        -- 'e'
        4 => (
        "00000000",
        "00000000",
        "00111000",
        "01000100",
        "01111000",
        "01000000",
        "00111000",
        "00000000"
        ),
        -- 'f'
        5 => (
        "00011000",
        "00100000",
        "01110000",
        "00100000",
        "00100000",
        "00100000",
        "00100000",
        "00000000"
        ),
        -- 'g'
        6 => (
        "00000000",
        "00111100",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'h'
        7 => (
        "01000000",
        "01000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00000000"
        ),
        -- 'i'
        8 => (
        "00010000",
        "00000000",
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- 'j'
        9 => (
        "00001000",
        "00000000",
        "00011000",
        "00001000",
        "00001000",
        "01001000",
        "00110000",
        "00000000"
        ),
        -- 'k'
        10 => (
        "01000000",
        "01010000",
        "01100000",
        "01110000",
        "01011000",
        "01001000",
        "01000100",
        "00000000"
        ),
        -- 'l'
        11 => (
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- 'm'
        12 => (
        "00000000",
        "00000000",
        "01101000",
        "01010100",
        "01010100",
        "01010100",
        "01010100",
        "00000000"
        ),
        -- 'n'
        13 => (
        "00000000",
        "00000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00000000"
        ),
        -- 'o'
        14 => (
        "00000000",
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- 'p'
        15 => (
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "01000000",
        "01000000",
        "00000000"
        ),
        -- 'q'
        16 => (
        "00000000",
        "00111100",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00000000"
        ),
        -- 'r'
        17 => (
        "00000000",
        "00000000",
        "01011000",
        "01100100",
        "01000000",
        "01000000",
        "01000000",
        "00000000"
        ),
        -- 's'
        18 => (
        "00000000",
        "00000000",
        "00111100",
        "01000000",
        "00111000",
        "00000100",
        "01111000",
        "00000000"
        ),
        -- 't'
        19 => (
        "00100000",
        "00100000",
        "01110000",
        "00100000",
        "00100000",
        "00100000",
        "00011000",
        "00000000"
        ),
        -- 'u'
        20 => (
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00111000",
        "00000000"
        ),
        -- 'v'
        21 => (
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "01001000",
        "00110000",
        "00010000",
        "00000000"
        ),
        -- 'w'
        22 => (
        "00000000",
        "00000000",
        "01000100",
        "01010100",
        "01010100",
        "01111100",
        "01000100",
        "00000000"
        ),
        -- 'x'
        23 => (
        "00000000",
        "00000000",
        "01000100",
        "00101000",
        "00010000",
        "00101000",
        "01000100",
        "00000000"
        ),
        -- 'y'
        24 => (
        "00000000",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'z'
        25 => (
        "00000000",
        "00000000",
        "01111100",
        "00001000",
        "00010000",
        "00100000",
        "01111100",
        "00000000"
        ),
        -- '0'
        26 => (
        "00111000",
        "01000100",
        "01001100",
        "01010100",
        "01100100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '1'
        27 => (
        "00010000",
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- '2'
        28 => (
        "00111000",
        "01000100",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "01111100",
        "00000000"
        ),
        -- '3'
        29 => (
        "00111000",
        "01000100",
        "00000100",
        "00011000",
        "00000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '4'
        30 => (
        "00001000",
        "00011000",
        "00101000",
        "01001000",
        "01111100",
        "00001000",
        "00001000",
        "00000000"
        ),
        -- '5'
        31 => (
        "01111100",
        "01000000",
        "01111000",
        "00000100",
        "00000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '6'
        32 => (
        "00111000",
        "01000000",
        "01000000",
        "01111000",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '7'
        33 => (
        "01111100",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "00100000",
        "00100000",
        "00000000"
        ),
        -- '8'
        34 => (
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '9'
        35 => (
        "00111000",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00111000",
        "00000000"
        )
    );
    signal index : integer;
begin
    index <= to_integer(unsigned(char_addr));

    -- Process to index into FONT_ROM using char_addr
    process (clk)
    begin
        if index < 36 then
            char_data <= FONT_ROM(index);
        else
            char_data <= (others => (others => '0'));
        end if;
    end process;

end rom;