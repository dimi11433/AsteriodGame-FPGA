library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Types.all;

entity get_character_rom is
    port (
        char_addr : in std_logic_vector(7 downto 0);
        char_data : out char_bitmap
    );
end entity get_character_rom;

architecture rom of get_character_rom is
    -- char_bitmap type is now declared in Font_Types package.
    -- Define a type for the complete font ROM: 26 letters + 10 digits = 36 characters.
    type font_rom_type is array (0 to 35) of char_bitmap;

    constant FONT_ROM : font_rom_type := (
        -- '0'
        0 => (
        "00111000",
        "01000100",
        "01001100",
        "01010100",
        "01100100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '1'
        1 => (
        "00010000",
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- '2'
        2 => (
        "00111000",
        "01000100",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "01111100",
        "00000000"
        ),
        -- '3'
        3 => (
        "00111000",
        "01000100",
        "00000100",
        "00011000",
        "00000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '4'
        4 => (
        "00001000",
        "00011000",
        "00101000",
        "01001000",
        "01111100",
        "00001000",
        "00001000",
        "00000000"
        ),
        -- '5'
        5 => (
        "01111100",
        "01000000",
        "01111000",
        "00000100",
        "00000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '6'
        6 => (
        "00111000",
        "01000000",
        "01000000",
        "01111000",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '7'
        7 => (
        "01111100",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "00100000",
        "00100000",
        "00000000"
        ),
        -- '8'
        8 => (
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- '9'
        9 => (
        "00111000",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'a'
        10 => (
        "00000000",
        "00000000",
        "00111000",
        "00000100",
        "00111100",
        "01000100",
        "00111100",
        "00000000"
        ),
        -- 'b'
        11 => (
        "01000000",
        "01000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01110000",
        "00000000"
        ),
        -- 'c'
        12 => (
        "00000000",
        "00000000",
        "00111000",
        "01000000",
        "01000000",
        "01000000",
        "00111000",
        "00000000"
        ),
        -- 'd'
        13 => (
        "00000100",
        "00000100",
        "00110100",
        "01001100",
        "01000100",
        "01000100",
        "00111100",
        "00000000"
        ),
        -- 'e'
        14 => (
        "00000000",
        "00000000",
        "00111000",
        "01000100",
        "01111000",
        "01000000",
        "00111000",
        "00000000"
        ),
        -- 'f'
        15 => (
        "00011000",
        "00100000",
        "01110000",
        "00100000",
        "00100000",
        "00100000",
        "00100000",
        "00000000"
        ),
        -- 'g'
        16 => (
        "00000000",
        "00111100",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'h'
        17 => (
        "01000000",
        "01000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00000000"
        ),
        -- 'i'
        18 => (
        "00010000",
        "00000000",
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- 'j'
        19 => (
        "00001000",
        "00000000",
        "00011000",
        "00001000",
        "00001000",
        "01001000",
        "00110000",
        "00000000"
        ),
        -- 'k'
        20 => (
        "01000000",
        "01010000",
        "01100000",
        "01110000",
        "01011000",
        "01001000",
        "01000100",
        "00000000"
        ),
        -- 'l'
        21 => (
        "00110000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00010000",
        "00111000",
        "00000000"
        ),
        -- 'm'
        22 => (
        "00000000",
        "00000000",
        "01101000",
        "01010100",
        "01010100",
        "01010100",
        "01010100",
        "00000000"
        ),
        -- 'n'
        23 => (
        "00000000",
        "00000000",
        "01110000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00000000"
        ),
        -- 'o'
        24 => (
        "00000000",
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "01000100",
        "00111000",
        "00000000"
        ),
        -- 'p'
        25 => (
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "00111000",
        "01000000",
        "01000000",
        "00000000"
        ),
        -- 'q'
        26 => (
        "00000000",
        "00111100",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00000000"
        ),
        -- 'r'
        27 => (
        "00000000",
        "00000000",
        "01011000",
        "01100100",
        "01000000",
        "01000000",
        "01000000",
        "00000000"
        ),
        -- 's'
        28 => (
        "00000000",
        "00000000",
        "00111100",
        "01000000",
        "00111000",
        "00000100",
        "01111000",
        "00000000"
        ),
        -- 't'
        29 => (
        "00100000",
        "00100000",
        "01110000",
        "00100000",
        "00100000",
        "00100000",
        "00011000",
        "00000000"
        ),
        -- 'u'
        30 => (
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "01001000",
        "01001000",
        "00111000",
        "00000000"
        ),
        -- 'v'
        31 => (
        "00000000",
        "00000000",
        "01001000",
        "01001000",
        "01001000",
        "00110000",
        "00010000",
        "00000000"
        ),
        -- 'w'
        32 => (
        "00000000",
        "00000000",
        "01000100",
        "01010100",
        "01010100",
        "01111100",
        "01000100",
        "00000000"
        ),
        -- 'x'
        33 => (
        "00000000",
        "00000000",
        "01000100",
        "00101000",
        "00010000",
        "00101000",
        "01000100",
        "00000000"
        ),
        -- 'y'
        34 => (
        "00000000",
        "01000100",
        "01000100",
        "00111100",
        "00000100",
        "00000100",
        "00111000",
        "00000000"
        ),
        -- 'z'
        35 => (
        "00000000",
        "00000000",
        "01111100",
        "00001000",
        "00010000",
        "00100000",
        "01111100",
        "00000000"
        )
    );
    signal index : integer;
begin
    index <= to_integer(unsigned(char_addr));

    -- Process to index into FONT_ROM using char_addr
    process (clk)
    begin
        if index < 36 then
            char_data <= FONT_ROM(index);
        else
            char_data <= (others => (others => '0'));
        end if;
    end process;

end rom;